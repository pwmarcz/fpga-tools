`include "uart_memory.v"

module Top;
  reg clock;
  reg received = 0;
  reg [7:0] rx_byte;

  wire transmit;
  wire [7:0] tx_byte;

  memory_controller mc(clock, received, rx_byte, transmit, tx_byte);

  initial
    begin
      $monitor($time,
               " clock = %d, received = %H, rx_byte = %H, transmit = %H, tx_byte = %H",
               clock, received, rx_byte, transmit, tx_byte);

      $dumpfile("controller_tb.vcd");
      $dumpvars;
    end

  initial
    begin
      clock = 0;
      forever #1 clock = ~clock;
    end

  task recv_byte;
    input [7:0] b;
    begin
      #2 received = 1; rx_byte = b;
      #2 received = 0;
    end
  endtask // recv_byte

  initial
    begin
      received = 0;

      recv_byte(`COMMAND_WRITE);
      recv_byte(3);
      recv_byte('h0E);
      recv_byte('hCD);
      recv_byte('h42);
      recv_byte('h43);
      recv_byte('h44);

      recv_byte(`COMMAND_WRITE);
      recv_byte(3);
      recv_byte('h0A);
      recv_byte('h10);
      recv_byte('h44);
      recv_byte('h45);
      recv_byte('h46);

      #2 recv_byte(`COMMAND_READ);
      recv_byte(1);
      recv_byte('h0E);
      recv_byte('hCD);

      #2 recv_byte(`COMMAND_READ);
      recv_byte(1);
      recv_byte('h0A);
      recv_byte('h10);

      #2 $finish;

    end

endmodule // Top
